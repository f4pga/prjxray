/*
ROM128X1: 128-Deep by 1-Wide ROM
ROM256X1: 256-Deep by 1-Wide ROM
ROM32X1: 32-Deep by 1-Wide ROM
ROM64X1: 64-Deep by 1-Wide ROM
*/

module top(input clk, stb, di, output do);
	localparam integer DIN_N = 256;
	localparam integer DOUT_N = 256;

	reg [DIN_N-1:0] din;
	wire [DOUT_N-1:0] dout;

	reg [DIN_N-1:0] din_shr;
	reg [DOUT_N-1:0] dout_shr;

	always @(posedge clk) begin
		din_shr <= {din_shr, di};
		dout_shr <= {dout_shr, din_shr[DIN_N-1]};
		if (stb) begin
			din <= din_shr;
			dout_shr <= dout;
		end
	end

	assign do = dout_shr[DOUT_N-1];

	roi roi (
		.clk(clk),
		.din(din),
		.dout(dout)
	);
endmodule

module roi(input clk, input [255:0] din, output [255:0] dout);
    ram_RAMB18E1 #(.LOC("XXX"))
            ram_RAMB18E1(.clk(clk), .din(din[  0 +: 8]), .dout(dout[  0 +: 8]));
endmodule

/*
Site RAMB18_X0Y42
Pushed it outside the pblock
lets extend pblock
*/
module ram_RAMB18E1 (input clk, input [7:0] din, output [7:0] dout);
    parameter LOC = "";

    RAMB18E1 #(
            .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .IS_CLKARDCLK_INVERTED(1'b0),
            .IS_CLKBWRCLK_INVERTED(1'b0),
            .IS_ENARDEN_INVERTED(1'b0),
            .IS_ENBWREN_INVERTED(1'b0),
            .IS_RSTRAMARSTRAM_INVERTED(1'b0),
            .IS_RSTRAMB_INVERTED(1'b0),
            .IS_RSTREGARSTREG_INVERTED(1'b0),
            .IS_RSTREGB_INVERTED(1'b0),
            .RAM_MODE("TDP"),
            .WRITE_MODE_A("WRITE_FIRST"),
            .WRITE_MODE_B("WRITE_FIRST"),
            .SIM_DEVICE("VIRTEX6")
        ) ram (
            .CLKARDCLK(din[0]),
            .CLKBWRCLK(din[1]),
            .ENARDEN(din[2]),
            .ENBWREN(din[3]),
            .REGCEAREGCE(din[4]),
            .REGCEB(din[5]),
            .RSTRAMARSTRAM(din[6]),
            .RSTRAMB(din[7]),
            .RSTREGARSTREG(din[0]),
            .RSTREGB(din[1]),
            .ADDRARDADDR(din[2]),
            .ADDRBWRADDR(din[3]),
            .DIADI(din[4]),
            .DIBDI(din[5]),
            .DIPADIP(din[6]),
            .DIPBDIP(din[7]),
            .WEA(din[0]),
            .WEBWE(din[1]),
            .DOADO(dout[0]),
            .DOBDO(dout[1]),
            .DOPADOP(dout[2]),
            .DOPBDOP(dout[3]));

endmodule

module ram_RAMB36E1 (input clk, input [7:0] din, output [7:0] dout);
    parameter LOC = "";

    RAMB36E1 #(
            .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            .IS_CLKARDCLK_INVERTED(1'b0),
            .IS_CLKBWRCLK_INVERTED(1'b0),
            .IS_ENARDEN_INVERTED(1'b0),
            .IS_ENBWREN_INVERTED(1'b0),
            .IS_RSTRAMARSTRAM_INVERTED(1'b0),
            .IS_RSTRAMB_INVERTED(1'b0),
            .IS_RSTREGARSTREG_INVERTED(1'b0),
            .IS_RSTREGB_INVERTED(1'b0),
            .RAM_MODE("TDP"),
            .WRITE_MODE_A("WRITE_FIRST"),
            .WRITE_MODE_B("WRITE_FIRST"),
            .SIM_DEVICE("VIRTEX6")
        ) ram (
            .CLKARDCLK(din[0]),
            .CLKBWRCLK(din[1]),
            .ENARDEN(din[2]),
            .ENBWREN(din[3]),
            .REGCEAREGCE(din[4]),
            .REGCEB(din[5]),
            .RSTRAMARSTRAM(din[6]),
            .RSTRAMB(din[7]),
            .RSTREGARSTREG(din[0]),
            .RSTREGB(din[1]),
            .ADDRARDADDR(din[2]),
            .ADDRBWRADDR(din[3]),
            .DIADI(din[4]),
            .DIBDI(din[5]),
            .DIPADIP(din[6]),
            .DIPBDIP(din[7]),
            .WEA(din[0]),
            .WEBWE(din[1]),
            .DOADO(dout[0]),
            .DOBDO(dout[1]),
            .DOPADOP(dout[2]),
            .DOPBDOP(dout[3]));
endmodule

