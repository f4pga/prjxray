module top(input di, output do);

   assign do = di;

endmodule
