
module top(input clk, ce, sr, d, output q);
	(* LOC="SLICE_X16Y100", BEL="AFF", DONT_TOUCH *)
	LDCE ff (
		.G(clk),
		.GE(ce),
		.CLR(sr),
		.D(d),
		.Q(q)
	);
endmodule

