`ifndef ROI
ERROR: must set ROI
`endif

module top(input clk, stb, di, output do);
	localparam integer DIN_N = 256;
	localparam integer DOUT_N = 256;

	reg [DIN_N-1:0] din;
	wire [DOUT_N-1:0] dout;

	reg [DIN_N-1:0] din_shr;
	reg [DOUT_N-1:0] dout_shr;

	always @(posedge clk) begin
		din_shr <= {din_shr, di};
		dout_shr <= {dout_shr, din_shr[DIN_N-1]};
		if (stb) begin
			din <= din_shr;
			dout_shr <= dout;
		end
	end

	assign do = dout_shr[DOUT_N-1];

    `ROI
	    roi (
		.clk(clk),
		.din(din),
		.dout(dout)
	);
endmodule

module roi_io_a(input clk, input [255:0] din, output [255:0] dout);
    assign dout[0] = din[0] & din[1];

    IOBUF_INTERMDISABLE #(
        .DRIVE(12),
        .IBUF_LOW_PWR("TRUE"),
        .IOSTANDARD("DEFAULT"),
        .SLEW("SLOW"),
        .USE_IBUFDISABLE("TRUE")
    ) IOBUF_INTERMDISABLE_inst (
        .O(1'b0),
        .IO(1'bz),
        .I(dout[8]),
        .IBUFDISABLE(1'b0),
        .INTERMDISABLE(1'b0),
        .T(1'b1));

endmodule

module roi_io_b(input clk, input [255:0] din, output [255:0] dout);
    assign dout[0] = din[0] & din[1];

    wire onet;

    IOBUF_INTERMDISABLE #(
        .DRIVE(12),
        .IBUF_LOW_PWR("FALSE"),
        .IOSTANDARD("DEFAULT"),
        .SLEW("SLOW"),
        .USE_IBUFDISABLE("FALSE")
    ) IOBUF_INTERMDISABLE_inst (
        .O(onet),
        .IO(1'bz),
        .I(dout[8]),
        .IBUFDISABLE(1'b0),
        .INTERMDISABLE(1'b0),
        .T(1'b1));

    PULLUP PULLUP_inst (
        .O(onet)
    );

    IOBUF_INTERMDISABLE #(
        .DRIVE(12),
        .IBUF_LOW_PWR("FALSE"),
        .IOSTANDARD("DEFAULT"),
        .SLEW("SLOW"),
        .USE_IBUFDISABLE("FALSE")
    ) i2 (
        .O(),
        .IO(1'bz),
        .I(dout[8]),
        .IBUFDISABLE(1'b0),
        .INTERMDISABLE(1'b0),
        .T(1'b1));

endmodule

