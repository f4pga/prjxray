module top (input a, b, c, output x, y, z);
	assign x = a, y = b, z = c;
endmodule
